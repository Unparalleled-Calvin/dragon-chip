`ifndef __MYCOMMON_SVH__
`define __MYCOMMON_SVH__

`include "common.svh"

typedef `BITS(10) i10;
typedef `BITS(20) i20;
typedef `BITS(22) i22;

`endif
